module hex_to_7seg (in0_3,in4_7,in8_9,out0_3,out4_7,out8_9);

	output [6:0] out0_3;
	input [3:0] in0_3;
	reg [6:0] out0_3;
	
	//same logic as 0-3
	output [6:0] out4_7;
	input [3:0] in4_7;
	reg [6:0] out4_7;
	
	output [6:0] out8_9;
	input [1:0] in8_9;
	reg [6:0] out8_9;
	
	always @ (*)
		case (in0_3)
			4'h0: out0_3 = 7'b1000000;
			4'h1: out0_3 = 7'b1111001;
			4'h2: out0_3 = 7'b0100100;
			4'h3: out0_3 = 7'b0110000;
			4'h4: out0_3 = 7'b0011001;
			4'h5: out0_3 = 7'b0010010;
			4'h6: out0_3 = 7'b0000010;
			4'h7: out0_3 = 7'b1111000;
			4'h8: out0_3 = 7'b0000000;
			4'h9: out0_3 = 7'b0011000;
			4'ha: out0_3 = 7'b0001000;
			4'hb: out0_3 = 7'b0000011;
			4'hc: out0_3 = 7'b1000110;
			4'hd: out0_3 = 7'b0100001;
			4'he: out0_3 = 7'b0000110;
			4'hf: out0_3 = 7'b0001110;
		endcase
	
	always @ (*)		
		case (in4_7)
			4'h0: out4_7 = 7'b1000000;
			4'h1: out4_7 = 7'b1111001;
			4'h2: out4_7 = 7'b0100100;
			4'h3: out4_7 = 7'b0110000;
			4'h4: out4_7 = 7'b0011001;
			4'h5: out4_7 = 7'b0010010;
			4'h6: out4_7 = 7'b0000010;
			4'h7: out4_7 = 7'b1111000;
			4'h8: out4_7 = 7'b0000000;
			4'h9: out4_7 = 7'b0011000;
			4'ha: out4_7 = 7'b0001000;
			4'hb: out4_7 = 7'b0000011;
			4'hc: out4_7 = 7'b1000110;
			4'hd: out4_7 = 7'b0100001;
			4'he: out4_7 = 7'b0000110;
			4'hf: out4_7 = 7'b0001110;
		endcase
	
	always @ (*)
		case (in8_9)
			4'h0: out8_9 = 7'b1000000;
			4'h1: out8_9 = 7'b1111001;
			4'h2: out8_9 = 7'b0100100;
			4'h3: out8_9 = 7'b0110000;
		endcase

endmodule
